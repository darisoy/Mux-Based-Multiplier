module cell1(input  logic xj, yj, sin, cin, xi, yi, si
             output logic cout, sout);

    logic temp0;
    4_1_mux    cell1_mux (.in0(1'b0), .in1(yi), .in2(xi), .in3(si), .sel0(xj), .sel1(yj), .out(temp0));
    full_adder cell1_fa  (.in0(temp0), .in1(sin), .cin(cin), .sum(sout), .cout(cout));

endmodule
